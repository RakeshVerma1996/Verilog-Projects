
module SR_FLIP(input wire S,
               input wire R,
               input wire clk,
               input wire reset,
         
  
